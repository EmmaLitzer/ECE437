
`timescale 1ns / 1ps

module FSM(    
    output [7:0] led,
    input  sys_clkn,
    input  sys_clkp,
    output ADT7420_A0,
    output ADT7420_A1,
    output I2C_SCL_0,
    inout  I2C_SDA_0,        
    output reg FSM_Clk_reg,    
    output reg ILA_Clk_reg,
    output reg ACK_bit,
    output reg SCL,
    output reg SDA,
    output reg [7:0] State,
    output wire [31:0] PCDATA,
    output wire [31:0] STARTR,
    output wire [31:0] STARTW,
    input  wire    [4:0] okUH,
    output wire    [2:0] okHU,
    inout  wire    [31:0] okUHU,   
    inout wire okAA     
    );
    
    
    //Instantiate the ClockGenerator module, where three signals are generate:
    //High speed CLK signal, Low speed FSM_Clk signal     
    wire [23:0] ClkDivThreshold = 100;   
    wire FSM_Clk, ILA_Clk; 
    ClockGenerator ClockGenerator1 (  .sys_clkn(sys_clkn),
                                      .sys_clkp(sys_clkp),                                      
                                      .ClkDivThreshold(ClkDivThreshold),
                                      .FSM_Clk(FSM_Clk),                                      
                                      .ILA_Clk(ILA_Clk) );
    
                                        
    wire [6:0] devaddrw = PCDATA[31:23];
    wire [6:0] devaddrr = PCDATA[15:7];
    wire [7:0] regaddr = PCDATA[23:16];
    wire RW = PCDATA[0]; //should always be 1
    wire currstate;
    wire error_bit;
    wire MSB;
    wire LSB;   
    
    Write write2read (  .devaddr(devaddrw),
                        .regaddr(regaddr),
                        .START(STARTW[0]),
                        .I2C_SCL_0(I2C_SCL_0),
                        .I2C_SDA_0(I2C_SDA_0),
                        .SCL(SCL),
                        .SDA(SDA),
                        .FSM_Clk(FSM_Clk),                                      
                        .ILA_Clk(ILA_Clk),
                        .ILA_Clk(ILA_Clk),
                        .FSM_Clk_reg(FSM_Clk_reg),
                        .ILA_Clk_reg(ILA_Clk_reg),
                        .State(currstate),
                        .ACK_bit(ACK_bit),
                        .error_bit(error_bit)
                      );
                      
    Read read_data (    .devaddr(devaddrr),
                        .DATAL(LSB),
                        .DATAH(MSB),
                        .START(STARTR[0]),
                        .I2C_SCL_0(I2C_SCL_0),
                        .I2C_SDA_0(I2C_SDA_0),
                        .SCL(SCL),
                        .SDA(SDA),
                        .FSM_Clk(FSM_Clk),                                      
                        .ILA_Clk(ILA_Clk),
                        .FSM_Clk_reg(FSM_Clk_reg),
                        .ILA_Clk_reg(ILA_Clk_reg),
                        .State(currstate),
                        .ACK_bit(ACK_bit),
                        .error_bit(error_bit)
                      );     
       
    localparam STATE_INIT       = 8'd0;    
    assign led[7] = ACK_bit;
    assign led[6] = error_bit;                         
    
    // OK Interface
    wire [112:0]    okHE;  //These are FrontPanel wires needed to IO communication    
    wire [64:0]     okEH;  //These are FrontPanel wires needed to IO communication 
        //Depending on the number of outgoing endpoints, adjust endPt_count accordingly.
    //In this example, we have 2 output endpoints, hence endPt_count = 2.
    localparam  endPt_count = 2;
    wire [endPt_count*65-1:0] okEHx;  
    okWireOR # (.N(endPt_count)) wireOR (okEH, okEHx);
    wire okClk;
    
    //This is the OK host that allows data to be sent or recived    
    okHost hostIF (
        .okUH(okUH),
        .okHU(okHU),
        .okUHU(okUHU),
        .okClk(okClk),
        .okAA(okAA),
        .okHE(okHE),
        .okEH(okEH)
    );
    
    //  PC_controll is a wire that contains data sent from the PC to FPGA.
    //  The data is communicated via memeory location 0x00
   okWireIn wire10 (   .okHE(okHE), 
                       .ep_addr(8'h00), 
                       .ep_dataout(PCDATA));  
                       
   okWireIn wire11 (   .okHE(okHE), 
                       .ep_addr(8'h01), 
                       .ep_dataout(STARTW));  
                       
    okWireIn wire12 (   .okHE(okHE), 
                       .ep_addr(8'h02), 
                       .ep_dataout(STARTR));                                                                                    
                      
   okWireOut wire21 (  .okHE(okHE), 
                   .okEH(okEHx[ 1*65 +: 65 ]), //unsure what this line is for but is giving errors
                   .ep_addr(8'h21), 
                   .ep_datain(MSB));
                  
   okWireOut wire20 (  .okHE(okHE), 
                   .okEH(okEHx[ 0*65 +: 65 ]),
                   .ep_addr(8'h20), 
                   .ep_datain(LSB));             
               
endmodule

`timescale 1ns / 1ps

module Testbench();
    //Declare wires and registers that will interface with the module under test
    //Registers are initilized to known states. Wires cannot be initilized.                 
    reg sys_clkn=1;
    wire sys_clkp;
    wire [7:0] led;
    reg [3:0] button;
    reg [31:0] PCDATA;
    wire [7:0] StateT;
    wire FSM_Clk_reg;
    reg [31:0] STARTW = 0;
    wire SDA;
    
    //Invoke the module that we like to test
    FSM ModuleUnderTest (.sys_clkn(sys_clkn), .sys_clkp(sys_clkp), .PCDATA(PCDATA), .State(StateT), .FSM_Clk_reg(FSM_Clk_reg), .STARTW(STARTW), .I2C_SDA_0(SDA));
    
    // Generate a clock signal. The clock will change its state every 5ns.
    //Remember that the test module takes sys_clkp and sys_clkn as input clock signals.
    //From these two signals a clock signal, clk, is derived.
    //The LVDS clock signal, sys_clkn, is always in the opposite state than sys_clkp.     
    assign sys_clkp = ~sys_clkn;    
    always begin
        #5 sys_clkn = ~sys_clkn;
    end        
      
    initial begin          
            #20000 PCDATA <= 32'b00110010001010000011001100000001;   
            #20000 STARTW <= 1;                                                   

            //#100 button <= 4'b1110;
          
    end

endmodule
